module test;



endmodule